`include "../tb/chaos_generator_tb.sv"
